
module sincos2 (
	clk,
	areset,
	a,
	c,
	s);	

	input		clk;
	input		areset;
	input	[9:0]	a;
	output	[4:0]	c;
	output	[4:0]	s;
endmodule

    Mac OS X            	   2   �      �                                      ATTR       �   �                     �     com.dropbox.attrs              com.dropbox.internal 

�s}�0^U�     ������
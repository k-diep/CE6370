// megafunction wizard: %RAM initializer%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTMEM_INIT 

// ============================================================
// File Name: ram1.v
// Megafunction Name(s):
// 			ALTMEM_INIT
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 22.1std.2 Build 922 07/20/2023 SC Lite Edition
// ************************************************************

//Copyright (C) 2023  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and any partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details, at
//https://fpgasoftware.intel.com/eula.

module ram1 (
	clock,
	init,
	dataout,
	init_busy,
	ram_address,
	ram_wren)/* synthesis synthesis_clearbox = 1 */;

	input	  clock;
	input	  init;
	output	[17:0]  dataout;
	output	  init_busy;
	output	[9:0]  ram_address;
	output	  ram_wren;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: INIT_FILE STRING "soc_system/syn/myproject_softmax_stable_ap_fixed_ap_fixed_16_6_5_3_0_softmax_config10_s_exp_table_ROM_bkb.mif"
// Retrieval info: CONSTANT: INIT_TO_ZERO STRING "NO"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altmem_init"
// Retrieval info: CONSTANT: NUMWORDS NUMERIC "1024"
// Retrieval info: CONSTANT: PORT_ROM_DATA_READY STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: ROM_READ_LATENCY NUMERIC "1"
// Retrieval info: CONSTANT: WIDTH NUMERIC "18"
// Retrieval info: CONSTANT: WIDTHAD NUMERIC "10"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: USED_PORT: dataout 0 0 18 0 OUTPUT NODEFVAL "dataout[17..0]"
// Retrieval info: CONNECT: dataout 0 0 18 0 @dataout 0 0 18 0
// Retrieval info: USED_PORT: init 0 0 0 0 INPUT NODEFVAL "init"
// Retrieval info: CONNECT: @init 0 0 0 0 init 0 0 0 0
// Retrieval info: USED_PORT: init_busy 0 0 0 0 OUTPUT NODEFVAL "init_busy"
// Retrieval info: CONNECT: init_busy 0 0 0 0 @init_busy 0 0 0 0
// Retrieval info: USED_PORT: ram_address 0 0 10 0 OUTPUT NODEFVAL "ram_address[9..0]"
// Retrieval info: CONNECT: ram_address 0 0 10 0 @ram_address 0 0 10 0
// Retrieval info: USED_PORT: ram_wren 0 0 0 0 OUTPUT NODEFVAL "ram_wren"
// Retrieval info: CONNECT: ram_wren 0 0 0 0 @ram_wren 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL ram1.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram1.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram1.bsf TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram1_inst.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram1_bb.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram1.inc TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram1.cmp TRUE TRUE
// Retrieval info: LIB_FILE: lpm
